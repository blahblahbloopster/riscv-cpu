0c_31d31b8d__00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_31d31b8d_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000
10_5cfbc662__00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_31d31b8d_00000000_00000000_00000000_5cfbc662_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000
10_e83c9fd7__00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_31d31b8d_00000000_00000000_00000000_e83c9fd7_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000
08_b7fc7fc0__00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_b7fc7fc0_00000000_00000000_00000000_31d31b8d_00000000_00000000_00000000_e83c9fd7_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000
1a_b616d702__00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_b7fc7fc0_00000000_00000000_00000000_31d31b8d_00000000_00000000_00000000_e83c9fd7_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_b616d702_00000000_00000000_00000000_00000000_00000000
19_d38b1ff2__00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_b7fc7fc0_00000000_00000000_00000000_31d31b8d_00000000_00000000_00000000_e83c9fd7_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_d38b1ff2_b616d702_00000000_00000000_00000000_00000000_00000000
1a_a3657290__00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_b7fc7fc0_00000000_00000000_00000000_31d31b8d_00000000_00000000_00000000_e83c9fd7_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_d38b1ff2_a3657290_00000000_00000000_00000000_00000000_00000000
06_07c6ecf4__00000000_00000000_00000000_00000000_00000000_00000000_07c6ecf4_00000000_b7fc7fc0_00000000_00000000_00000000_31d31b8d_00000000_00000000_00000000_e83c9fd7_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_d38b1ff2_a3657290_00000000_00000000_00000000_00000000_00000000
19_452a78ba__00000000_00000000_00000000_00000000_00000000_00000000_07c6ecf4_00000000_b7fc7fc0_00000000_00000000_00000000_31d31b8d_00000000_00000000_00000000_e83c9fd7_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_452a78ba_a3657290_00000000_00000000_00000000_00000000_00000000
09_eb3a9aa9__00000000_00000000_00000000_00000000_00000000_00000000_07c6ecf4_00000000_b7fc7fc0_eb3a9aa9_00000000_00000000_31d31b8d_00000000_00000000_00000000_e83c9fd7_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_452a78ba_a3657290_00000000_00000000_00000000_00000000_00000000
01_18aedfb7__00000000_18aedfb7_00000000_00000000_00000000_00000000_07c6ecf4_00000000_b7fc7fc0_eb3a9aa9_00000000_00000000_31d31b8d_00000000_00000000_00000000_e83c9fd7_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_452a78ba_a3657290_00000000_00000000_00000000_00000000_00000000
16_09b585e5__00000000_18aedfb7_00000000_00000000_00000000_00000000_07c6ecf4_00000000_b7fc7fc0_eb3a9aa9_00000000_00000000_31d31b8d_00000000_00000000_00000000_e83c9fd7_00000000_00000000_00000000_00000000_00000000_09b585e5_00000000_00000000_452a78ba_a3657290_00000000_00000000_00000000_00000000_00000000
1d_ba0054f6__00000000_18aedfb7_00000000_00000000_00000000_00000000_07c6ecf4_00000000_b7fc7fc0_eb3a9aa9_00000000_00000000_31d31b8d_00000000_00000000_00000000_e83c9fd7_00000000_00000000_00000000_00000000_00000000_09b585e5_00000000_00000000_452a78ba_a3657290_00000000_00000000_ba0054f6_00000000_00000000
14_53bfd2eb__00000000_18aedfb7_00000000_00000000_00000000_00000000_07c6ecf4_00000000_b7fc7fc0_eb3a9aa9_00000000_00000000_31d31b8d_00000000_00000000_00000000_e83c9fd7_00000000_00000000_00000000_53bfd2eb_00000000_09b585e5_00000000_00000000_452a78ba_a3657290_00000000_00000000_ba0054f6_00000000_00000000
19_0d056ce8__00000000_18aedfb7_00000000_00000000_00000000_00000000_07c6ecf4_00000000_b7fc7fc0_eb3a9aa9_00000000_00000000_31d31b8d_00000000_00000000_00000000_e83c9fd7_00000000_00000000_00000000_53bfd2eb_00000000_09b585e5_00000000_00000000_0d056ce8_a3657290_00000000_00000000_ba0054f6_00000000_00000000
0a_dee912e6__00000000_18aedfb7_00000000_00000000_00000000_00000000_07c6ecf4_00000000_b7fc7fc0_eb3a9aa9_dee912e6_00000000_31d31b8d_00000000_00000000_00000000_e83c9fd7_00000000_00000000_00000000_53bfd2eb_00000000_09b585e5_00000000_00000000_0d056ce8_a3657290_00000000_00000000_ba0054f6_00000000_00000000
04_b093df3b__00000000_18aedfb7_00000000_00000000_b093df3b_00000000_07c6ecf4_00000000_b7fc7fc0_eb3a9aa9_dee912e6_00000000_31d31b8d_00000000_00000000_00000000_e83c9fd7_00000000_00000000_00000000_53bfd2eb_00000000_09b585e5_00000000_00000000_0d056ce8_a3657290_00000000_00000000_ba0054f6_00000000_00000000
01_92c5c34e__00000000_92c5c34e_00000000_00000000_b093df3b_00000000_07c6ecf4_00000000_b7fc7fc0_eb3a9aa9_dee912e6_00000000_31d31b8d_00000000_00000000_00000000_e83c9fd7_00000000_00000000_00000000_53bfd2eb_00000000_09b585e5_00000000_00000000_0d056ce8_a3657290_00000000_00000000_ba0054f6_00000000_00000000
11_0eee3f38__00000000_92c5c34e_00000000_00000000_b093df3b_00000000_07c6ecf4_00000000_b7fc7fc0_eb3a9aa9_dee912e6_00000000_31d31b8d_00000000_00000000_00000000_e83c9fd7_0eee3f38_00000000_00000000_53bfd2eb_00000000_09b585e5_00000000_00000000_0d056ce8_a3657290_00000000_00000000_ba0054f6_00000000_00000000
0f_84d92790__00000000_92c5c34e_00000000_00000000_b093df3b_00000000_07c6ecf4_00000000_b7fc7fc0_eb3a9aa9_dee912e6_00000000_31d31b8d_00000000_00000000_84d92790_e83c9fd7_0eee3f38_00000000_00000000_53bfd2eb_00000000_09b585e5_00000000_00000000_0d056ce8_a3657290_00000000_00000000_ba0054f6_00000000_00000000
1e_393cfdf9__00000000_92c5c34e_00000000_00000000_b093df3b_00000000_07c6ecf4_00000000_b7fc7fc0_eb3a9aa9_dee912e6_00000000_31d31b8d_00000000_00000000_84d92790_e83c9fd7_0eee3f38_00000000_00000000_53bfd2eb_00000000_09b585e5_00000000_00000000_0d056ce8_a3657290_00000000_00000000_ba0054f6_393cfdf9_00000000
18_2cf5a75f__00000000_92c5c34e_00000000_00000000_b093df3b_00000000_07c6ecf4_00000000_b7fc7fc0_eb3a9aa9_dee912e6_00000000_31d31b8d_00000000_00000000_84d92790_e83c9fd7_0eee3f38_00000000_00000000_53bfd2eb_00000000_09b585e5_00000000_2cf5a75f_0d056ce8_a3657290_00000000_00000000_ba0054f6_393cfdf9_00000000
07_041ba92d__00000000_92c5c34e_00000000_00000000_b093df3b_00000000_07c6ecf4_041ba92d_b7fc7fc0_eb3a9aa9_dee912e6_00000000_31d31b8d_00000000_00000000_84d92790_e83c9fd7_0eee3f38_00000000_00000000_53bfd2eb_00000000_09b585e5_00000000_2cf5a75f_0d056ce8_a3657290_00000000_00000000_ba0054f6_393cfdf9_00000000
02_7b16b023__00000000_92c5c34e_7b16b023_00000000_b093df3b_00000000_07c6ecf4_041ba92d_b7fc7fc0_eb3a9aa9_dee912e6_00000000_31d31b8d_00000000_00000000_84d92790_e83c9fd7_0eee3f38_00000000_00000000_53bfd2eb_00000000_09b585e5_00000000_2cf5a75f_0d056ce8_a3657290_00000000_00000000_ba0054f6_393cfdf9_00000000
16_da967749__00000000_92c5c34e_7b16b023_00000000_b093df3b_00000000_07c6ecf4_041ba92d_b7fc7fc0_eb3a9aa9_dee912e6_00000000_31d31b8d_00000000_00000000_84d92790_e83c9fd7_0eee3f38_00000000_00000000_53bfd2eb_00000000_da967749_00000000_2cf5a75f_0d056ce8_a3657290_00000000_00000000_ba0054f6_393cfdf9_00000000
0a_88907a80__00000000_92c5c34e_7b16b023_00000000_b093df3b_00000000_07c6ecf4_041ba92d_b7fc7fc0_eb3a9aa9_88907a80_00000000_31d31b8d_00000000_00000000_84d92790_e83c9fd7_0eee3f38_00000000_00000000_53bfd2eb_00000000_da967749_00000000_2cf5a75f_0d056ce8_a3657290_00000000_00000000_ba0054f6_393cfdf9_00000000
00_e4cdda62__00000000_92c5c34e_7b16b023_00000000_b093df3b_00000000_07c6ecf4_041ba92d_b7fc7fc0_eb3a9aa9_88907a80_00000000_31d31b8d_00000000_00000000_84d92790_e83c9fd7_0eee3f38_00000000_00000000_53bfd2eb_00000000_da967749_00000000_2cf5a75f_0d056ce8_a3657290_00000000_00000000_ba0054f6_393cfdf9_00000000
1d_6eb08e55__00000000_92c5c34e_7b16b023_00000000_b093df3b_00000000_07c6ecf4_041ba92d_b7fc7fc0_eb3a9aa9_88907a80_00000000_31d31b8d_00000000_00000000_84d92790_e83c9fd7_0eee3f38_00000000_00000000_53bfd2eb_00000000_da967749_00000000_2cf5a75f_0d056ce8_a3657290_00000000_00000000_6eb08e55_393cfdf9_00000000
0c_4646d520__00000000_92c5c34e_7b16b023_00000000_b093df3b_00000000_07c6ecf4_041ba92d_b7fc7fc0_eb3a9aa9_88907a80_00000000_4646d520_00000000_00000000_84d92790_e83c9fd7_0eee3f38_00000000_00000000_53bfd2eb_00000000_da967749_00000000_2cf5a75f_0d056ce8_a3657290_00000000_00000000_6eb08e55_393cfdf9_00000000
05_e4c5244e__00000000_92c5c34e_7b16b023_00000000_b093df3b_e4c5244e_07c6ecf4_041ba92d_b7fc7fc0_eb3a9aa9_88907a80_00000000_4646d520_00000000_00000000_84d92790_e83c9fd7_0eee3f38_00000000_00000000_53bfd2eb_00000000_da967749_00000000_2cf5a75f_0d056ce8_a3657290_00000000_00000000_6eb08e55_393cfdf9_00000000
13_17906fda__00000000_92c5c34e_7b16b023_00000000_b093df3b_e4c5244e_07c6ecf4_041ba92d_b7fc7fc0_eb3a9aa9_88907a80_00000000_4646d520_00000000_00000000_84d92790_e83c9fd7_0eee3f38_00000000_17906fda_53bfd2eb_00000000_da967749_00000000_2cf5a75f_0d056ce8_a3657290_00000000_00000000_6eb08e55_393cfdf9_00000000
15_e468951c__00000000_92c5c34e_7b16b023_00000000_b093df3b_e4c5244e_07c6ecf4_041ba92d_b7fc7fc0_eb3a9aa9_88907a80_00000000_4646d520_00000000_00000000_84d92790_e83c9fd7_0eee3f38_00000000_17906fda_53bfd2eb_e468951c_da967749_00000000_2cf5a75f_0d056ce8_a3657290_00000000_00000000_6eb08e55_393cfdf9_00000000
16_52e30da7__00000000_92c5c34e_7b16b023_00000000_b093df3b_e4c5244e_07c6ecf4_041ba92d_b7fc7fc0_eb3a9aa9_88907a80_00000000_4646d520_00000000_00000000_84d92790_e83c9fd7_0eee3f38_00000000_17906fda_53bfd2eb_e468951c_52e30da7_00000000_2cf5a75f_0d056ce8_a3657290_00000000_00000000_6eb08e55_393cfdf9_00000000
1a_c72cb5ab__00000000_92c5c34e_7b16b023_00000000_b093df3b_e4c5244e_07c6ecf4_041ba92d_b7fc7fc0_eb3a9aa9_88907a80_00000000_4646d520_00000000_00000000_84d92790_e83c9fd7_0eee3f38_00000000_17906fda_53bfd2eb_e468951c_52e30da7_00000000_2cf5a75f_0d056ce8_c72cb5ab_00000000_00000000_6eb08e55_393cfdf9_00000000
0d_27348e13__00000000_92c5c34e_7b16b023_00000000_b093df3b_e4c5244e_07c6ecf4_041ba92d_b7fc7fc0_eb3a9aa9_88907a80_00000000_4646d520_27348e13_00000000_84d92790_e83c9fd7_0eee3f38_00000000_17906fda_53bfd2eb_e468951c_52e30da7_00000000_2cf5a75f_0d056ce8_c72cb5ab_00000000_00000000_6eb08e55_393cfdf9_00000000
06_9f459a20__00000000_92c5c34e_7b16b023_00000000_b093df3b_e4c5244e_9f459a20_041ba92d_b7fc7fc0_eb3a9aa9_88907a80_00000000_4646d520_27348e13_00000000_84d92790_e83c9fd7_0eee3f38_00000000_17906fda_53bfd2eb_e468951c_52e30da7_00000000_2cf5a75f_0d056ce8_c72cb5ab_00000000_00000000_6eb08e55_393cfdf9_00000000
10_c281ef89__00000000_92c5c34e_7b16b023_00000000_b093df3b_e4c5244e_9f459a20_041ba92d_b7fc7fc0_eb3a9aa9_88907a80_00000000_4646d520_27348e13_00000000_84d92790_c281ef89_0eee3f38_00000000_17906fda_53bfd2eb_e468951c_52e30da7_00000000_2cf5a75f_0d056ce8_c72cb5ab_00000000_00000000_6eb08e55_393cfdf9_00000000
0c_fbd237fa__00000000_92c5c34e_7b16b023_00000000_b093df3b_e4c5244e_9f459a20_041ba92d_b7fc7fc0_eb3a9aa9_88907a80_00000000_fbd237fa_27348e13_00000000_84d92790_c281ef89_0eee3f38_00000000_17906fda_53bfd2eb_e468951c_52e30da7_00000000_2cf5a75f_0d056ce8_c72cb5ab_00000000_00000000_6eb08e55_393cfdf9_00000000
0a_30cfaebf__00000000_92c5c34e_7b16b023_00000000_b093df3b_e4c5244e_9f459a20_041ba92d_b7fc7fc0_eb3a9aa9_30cfaebf_00000000_fbd237fa_27348e13_00000000_84d92790_c281ef89_0eee3f38_00000000_17906fda_53bfd2eb_e468951c_52e30da7_00000000_2cf5a75f_0d056ce8_c72cb5ab_00000000_00000000_6eb08e55_393cfdf9_00000000
12_a9c44efc__00000000_92c5c34e_7b16b023_00000000_b093df3b_e4c5244e_9f459a20_041ba92d_b7fc7fc0_eb3a9aa9_30cfaebf_00000000_fbd237fa_27348e13_00000000_84d92790_c281ef89_0eee3f38_a9c44efc_17906fda_53bfd2eb_e468951c_52e30da7_00000000_2cf5a75f_0d056ce8_c72cb5ab_00000000_00000000_6eb08e55_393cfdf9_00000000
00_78c53ae0__00000000_92c5c34e_7b16b023_00000000_b093df3b_e4c5244e_9f459a20_041ba92d_b7fc7fc0_eb3a9aa9_30cfaebf_00000000_fbd237fa_27348e13_00000000_84d92790_c281ef89_0eee3f38_a9c44efc_17906fda_53bfd2eb_e468951c_52e30da7_00000000_2cf5a75f_0d056ce8_c72cb5ab_00000000_00000000_6eb08e55_393cfdf9_00000000
02_693868f3__00000000_92c5c34e_693868f3_00000000_b093df3b_e4c5244e_9f459a20_041ba92d_b7fc7fc0_eb3a9aa9_30cfaebf_00000000_fbd237fa_27348e13_00000000_84d92790_c281ef89_0eee3f38_a9c44efc_17906fda_53bfd2eb_e468951c_52e30da7_00000000_2cf5a75f_0d056ce8_c72cb5ab_00000000_00000000_6eb08e55_393cfdf9_00000000
07_8d8d5c0b__00000000_92c5c34e_693868f3_00000000_b093df3b_e4c5244e_9f459a20_8d8d5c0b_b7fc7fc0_eb3a9aa9_30cfaebf_00000000_fbd237fa_27348e13_00000000_84d92790_c281ef89_0eee3f38_a9c44efc_17906fda_53bfd2eb_e468951c_52e30da7_00000000_2cf5a75f_0d056ce8_c72cb5ab_00000000_00000000_6eb08e55_393cfdf9_00000000
16_378472ee__00000000_92c5c34e_693868f3_00000000_b093df3b_e4c5244e_9f459a20_8d8d5c0b_b7fc7fc0_eb3a9aa9_30cfaebf_00000000_fbd237fa_27348e13_00000000_84d92790_c281ef89_0eee3f38_a9c44efc_17906fda_53bfd2eb_e468951c_378472ee_00000000_2cf5a75f_0d056ce8_c72cb5ab_00000000_00000000_6eb08e55_393cfdf9_00000000
1f_8958a65f__00000000_92c5c34e_693868f3_00000000_b093df3b_e4c5244e_9f459a20_8d8d5c0b_b7fc7fc0_eb3a9aa9_30cfaebf_00000000_fbd237fa_27348e13_00000000_84d92790_c281ef89_0eee3f38_a9c44efc_17906fda_53bfd2eb_e468951c_378472ee_00000000_2cf5a75f_0d056ce8_c72cb5ab_00000000_00000000_6eb08e55_393cfdf9_8958a65f
03_ae445cca__00000000_92c5c34e_693868f3_ae445cca_b093df3b_e4c5244e_9f459a20_8d8d5c0b_b7fc7fc0_eb3a9aa9_30cfaebf_00000000_fbd237fa_27348e13_00000000_84d92790_c281ef89_0eee3f38_a9c44efc_17906fda_53bfd2eb_e468951c_378472ee_00000000_2cf5a75f_0d056ce8_c72cb5ab_00000000_00000000_6eb08e55_393cfdf9_8958a65f
0b_de45cf71__00000000_92c5c34e_693868f3_ae445cca_b093df3b_e4c5244e_9f459a20_8d8d5c0b_b7fc7fc0_eb3a9aa9_30cfaebf_de45cf71_fbd237fa_27348e13_00000000_84d92790_c281ef89_0eee3f38_a9c44efc_17906fda_53bfd2eb_e468951c_378472ee_00000000_2cf5a75f_0d056ce8_c72cb5ab_00000000_00000000_6eb08e55_393cfdf9_8958a65f
01_0e710e6d__00000000_0e710e6d_693868f3_ae445cca_b093df3b_e4c5244e_9f459a20_8d8d5c0b_b7fc7fc0_eb3a9aa9_30cfaebf_de45cf71_fbd237fa_27348e13_00000000_84d92790_c281ef89_0eee3f38_a9c44efc_17906fda_53bfd2eb_e468951c_378472ee_00000000_2cf5a75f_0d056ce8_c72cb5ab_00000000_00000000_6eb08e55_393cfdf9_8958a65f
00_e1a0540a__00000000_0e710e6d_693868f3_ae445cca_b093df3b_e4c5244e_9f459a20_8d8d5c0b_b7fc7fc0_eb3a9aa9_30cfaebf_de45cf71_fbd237fa_27348e13_00000000_84d92790_c281ef89_0eee3f38_a9c44efc_17906fda_53bfd2eb_e468951c_378472ee_00000000_2cf5a75f_0d056ce8_c72cb5ab_00000000_00000000_6eb08e55_393cfdf9_8958a65f
15_da3000d4__00000000_0e710e6d_693868f3_ae445cca_b093df3b_e4c5244e_9f459a20_8d8d5c0b_b7fc7fc0_eb3a9aa9_30cfaebf_de45cf71_fbd237fa_27348e13_00000000_84d92790_c281ef89_0eee3f38_a9c44efc_17906fda_53bfd2eb_da3000d4_378472ee_00000000_2cf5a75f_0d056ce8_c72cb5ab_00000000_00000000_6eb08e55_393cfdf9_8958a65f
0b_ee7ca9a7__00000000_0e710e6d_693868f3_ae445cca_b093df3b_e4c5244e_9f459a20_8d8d5c0b_b7fc7fc0_eb3a9aa9_30cfaebf_ee7ca9a7_fbd237fa_27348e13_00000000_84d92790_c281ef89_0eee3f38_a9c44efc_17906fda_53bfd2eb_da3000d4_378472ee_00000000_2cf5a75f_0d056ce8_c72cb5ab_00000000_00000000_6eb08e55_393cfdf9_8958a65f
1d_4b162443__00000000_0e710e6d_693868f3_ae445cca_b093df3b_e4c5244e_9f459a20_8d8d5c0b_b7fc7fc0_eb3a9aa9_30cfaebf_ee7ca9a7_fbd237fa_27348e13_00000000_84d92790_c281ef89_0eee3f38_a9c44efc_17906fda_53bfd2eb_da3000d4_378472ee_00000000_2cf5a75f_0d056ce8_c72cb5ab_00000000_00000000_4b162443_393cfdf9_8958a65f
15_8042c02d__00000000_0e710e6d_693868f3_ae445cca_b093df3b_e4c5244e_9f459a20_8d8d5c0b_b7fc7fc0_eb3a9aa9_30cfaebf_ee7ca9a7_fbd237fa_27348e13_00000000_84d92790_c281ef89_0eee3f38_a9c44efc_17906fda_53bfd2eb_8042c02d_378472ee_00000000_2cf5a75f_0d056ce8_c72cb5ab_00000000_00000000_4b162443_393cfdf9_8958a65f
0f_05fb991e__00000000_0e710e6d_693868f3_ae445cca_b093df3b_e4c5244e_9f459a20_8d8d5c0b_b7fc7fc0_eb3a9aa9_30cfaebf_ee7ca9a7_fbd237fa_27348e13_00000000_05fb991e_c281ef89_0eee3f38_a9c44efc_17906fda_53bfd2eb_8042c02d_378472ee_00000000_2cf5a75f_0d056ce8_c72cb5ab_00000000_00000000_4b162443_393cfdf9_8958a65f
13_6282990b__00000000_0e710e6d_693868f3_ae445cca_b093df3b_e4c5244e_9f459a20_8d8d5c0b_b7fc7fc0_eb3a9aa9_30cfaebf_ee7ca9a7_fbd237fa_27348e13_00000000_05fb991e_c281ef89_0eee3f38_a9c44efc_6282990b_53bfd2eb_8042c02d_378472ee_00000000_2cf5a75f_0d056ce8_c72cb5ab_00000000_00000000_4b162443_393cfdf9_8958a65f
1e_1e097c79__00000000_0e710e6d_693868f3_ae445cca_b093df3b_e4c5244e_9f459a20_8d8d5c0b_b7fc7fc0_eb3a9aa9_30cfaebf_ee7ca9a7_fbd237fa_27348e13_00000000_05fb991e_c281ef89_0eee3f38_a9c44efc_6282990b_53bfd2eb_8042c02d_378472ee_00000000_2cf5a75f_0d056ce8_c72cb5ab_00000000_00000000_4b162443_1e097c79_8958a65f
12_d792537a__00000000_0e710e6d_693868f3_ae445cca_b093df3b_e4c5244e_9f459a20_8d8d5c0b_b7fc7fc0_eb3a9aa9_30cfaebf_ee7ca9a7_fbd237fa_27348e13_00000000_05fb991e_c281ef89_0eee3f38_d792537a_6282990b_53bfd2eb_8042c02d_378472ee_00000000_2cf5a75f_0d056ce8_c72cb5ab_00000000_00000000_4b162443_1e097c79_8958a65f
09_0683ab57__00000000_0e710e6d_693868f3_ae445cca_b093df3b_e4c5244e_9f459a20_8d8d5c0b_b7fc7fc0_0683ab57_30cfaebf_ee7ca9a7_fbd237fa_27348e13_00000000_05fb991e_c281ef89_0eee3f38_d792537a_6282990b_53bfd2eb_8042c02d_378472ee_00000000_2cf5a75f_0d056ce8_c72cb5ab_00000000_00000000_4b162443_1e097c79_8958a65f
0d_687d202e__00000000_0e710e6d_693868f3_ae445cca_b093df3b_e4c5244e_9f459a20_8d8d5c0b_b7fc7fc0_0683ab57_30cfaebf_ee7ca9a7_fbd237fa_687d202e_00000000_05fb991e_c281ef89_0eee3f38_d792537a_6282990b_53bfd2eb_8042c02d_378472ee_00000000_2cf5a75f_0d056ce8_c72cb5ab_00000000_00000000_4b162443_1e097c79_8958a65f
00_66f04107__00000000_0e710e6d_693868f3_ae445cca_b093df3b_e4c5244e_9f459a20_8d8d5c0b_b7fc7fc0_0683ab57_30cfaebf_ee7ca9a7_fbd237fa_687d202e_00000000_05fb991e_c281ef89_0eee3f38_d792537a_6282990b_53bfd2eb_8042c02d_378472ee_00000000_2cf5a75f_0d056ce8_c72cb5ab_00000000_00000000_4b162443_1e097c79_8958a65f
11_974251c3__00000000_0e710e6d_693868f3_ae445cca_b093df3b_e4c5244e_9f459a20_8d8d5c0b_b7fc7fc0_0683ab57_30cfaebf_ee7ca9a7_fbd237fa_687d202e_00000000_05fb991e_c281ef89_974251c3_d792537a_6282990b_53bfd2eb_8042c02d_378472ee_00000000_2cf5a75f_0d056ce8_c72cb5ab_00000000_00000000_4b162443_1e097c79_8958a65f
01_95aefe44__00000000_95aefe44_693868f3_ae445cca_b093df3b_e4c5244e_9f459a20_8d8d5c0b_b7fc7fc0_0683ab57_30cfaebf_ee7ca9a7_fbd237fa_687d202e_00000000_05fb991e_c281ef89_974251c3_d792537a_6282990b_53bfd2eb_8042c02d_378472ee_00000000_2cf5a75f_0d056ce8_c72cb5ab_00000000_00000000_4b162443_1e097c79_8958a65f
0e_d3095e51__00000000_95aefe44_693868f3_ae445cca_b093df3b_e4c5244e_9f459a20_8d8d5c0b_b7fc7fc0_0683ab57_30cfaebf_ee7ca9a7_fbd237fa_687d202e_d3095e51_05fb991e_c281ef89_974251c3_d792537a_6282990b_53bfd2eb_8042c02d_378472ee_00000000_2cf5a75f_0d056ce8_c72cb5ab_00000000_00000000_4b162443_1e097c79_8958a65f
10_76f15d5d__00000000_95aefe44_693868f3_ae445cca_b093df3b_e4c5244e_9f459a20_8d8d5c0b_b7fc7fc0_0683ab57_30cfaebf_ee7ca9a7_fbd237fa_687d202e_d3095e51_05fb991e_76f15d5d_974251c3_d792537a_6282990b_53bfd2eb_8042c02d_378472ee_00000000_2cf5a75f_0d056ce8_c72cb5ab_00000000_00000000_4b162443_1e097c79_8958a65f
17_e66ba7c1__00000000_95aefe44_693868f3_ae445cca_b093df3b_e4c5244e_9f459a20_8d8d5c0b_b7fc7fc0_0683ab57_30cfaebf_ee7ca9a7_fbd237fa_687d202e_d3095e51_05fb991e_76f15d5d_974251c3_d792537a_6282990b_53bfd2eb_8042c02d_378472ee_e66ba7c1_2cf5a75f_0d056ce8_c72cb5ab_00000000_00000000_4b162443_1e097c79_8958a65f
15_9bda402f__00000000_95aefe44_693868f3_ae445cca_b093df3b_e4c5244e_9f459a20_8d8d5c0b_b7fc7fc0_0683ab57_30cfaebf_ee7ca9a7_fbd237fa_687d202e_d3095e51_05fb991e_76f15d5d_974251c3_d792537a_6282990b_53bfd2eb_9bda402f_378472ee_e66ba7c1_2cf5a75f_0d056ce8_c72cb5ab_00000000_00000000_4b162443_1e097c79_8958a65f
15_4d24c9a9__00000000_95aefe44_693868f3_ae445cca_b093df3b_e4c5244e_9f459a20_8d8d5c0b_b7fc7fc0_0683ab57_30cfaebf_ee7ca9a7_fbd237fa_687d202e_d3095e51_05fb991e_76f15d5d_974251c3_d792537a_6282990b_53bfd2eb_4d24c9a9_378472ee_e66ba7c1_2cf5a75f_0d056ce8_c72cb5ab_00000000_00000000_4b162443_1e097c79_8958a65f
12_f9ea64b0__00000000_95aefe44_693868f3_ae445cca_b093df3b_e4c5244e_9f459a20_8d8d5c0b_b7fc7fc0_0683ab57_30cfaebf_ee7ca9a7_fbd237fa_687d202e_d3095e51_05fb991e_76f15d5d_974251c3_f9ea64b0_6282990b_53bfd2eb_4d24c9a9_378472ee_e66ba7c1_2cf5a75f_0d056ce8_c72cb5ab_00000000_00000000_4b162443_1e097c79_8958a65f
0d_2a7b62da__00000000_95aefe44_693868f3_ae445cca_b093df3b_e4c5244e_9f459a20_8d8d5c0b_b7fc7fc0_0683ab57_30cfaebf_ee7ca9a7_fbd237fa_2a7b62da_d3095e51_05fb991e_76f15d5d_974251c3_f9ea64b0_6282990b_53bfd2eb_4d24c9a9_378472ee_e66ba7c1_2cf5a75f_0d056ce8_c72cb5ab_00000000_00000000_4b162443_1e097c79_8958a65f
0e_1fdf13ab__00000000_95aefe44_693868f3_ae445cca_b093df3b_e4c5244e_9f459a20_8d8d5c0b_b7fc7fc0_0683ab57_30cfaebf_ee7ca9a7_fbd237fa_2a7b62da_1fdf13ab_05fb991e_76f15d5d_974251c3_f9ea64b0_6282990b_53bfd2eb_4d24c9a9_378472ee_e66ba7c1_2cf5a75f_0d056ce8_c72cb5ab_00000000_00000000_4b162443_1e097c79_8958a65f
0a_33a4289e__00000000_95aefe44_693868f3_ae445cca_b093df3b_e4c5244e_9f459a20_8d8d5c0b_b7fc7fc0_0683ab57_33a4289e_ee7ca9a7_fbd237fa_2a7b62da_1fdf13ab_05fb991e_76f15d5d_974251c3_f9ea64b0_6282990b_53bfd2eb_4d24c9a9_378472ee_e66ba7c1_2cf5a75f_0d056ce8_c72cb5ab_00000000_00000000_4b162443_1e097c79_8958a65f
18_46e91766__00000000_95aefe44_693868f3_ae445cca_b093df3b_e4c5244e_9f459a20_8d8d5c0b_b7fc7fc0_0683ab57_33a4289e_ee7ca9a7_fbd237fa_2a7b62da_1fdf13ab_05fb991e_76f15d5d_974251c3_f9ea64b0_6282990b_53bfd2eb_4d24c9a9_378472ee_e66ba7c1_46e91766_0d056ce8_c72cb5ab_00000000_00000000_4b162443_1e097c79_8958a65f
12_a22c7cf8__00000000_95aefe44_693868f3_ae445cca_b093df3b_e4c5244e_9f459a20_8d8d5c0b_b7fc7fc0_0683ab57_33a4289e_ee7ca9a7_fbd237fa_2a7b62da_1fdf13ab_05fb991e_76f15d5d_974251c3_a22c7cf8_6282990b_53bfd2eb_4d24c9a9_378472ee_e66ba7c1_46e91766_0d056ce8_c72cb5ab_00000000_00000000_4b162443_1e097c79_8958a65f
14_50f6b395__00000000_95aefe44_693868f3_ae445cca_b093df3b_e4c5244e_9f459a20_8d8d5c0b_b7fc7fc0_0683ab57_33a4289e_ee7ca9a7_fbd237fa_2a7b62da_1fdf13ab_05fb991e_76f15d5d_974251c3_a22c7cf8_6282990b_50f6b395_4d24c9a9_378472ee_e66ba7c1_46e91766_0d056ce8_c72cb5ab_00000000_00000000_4b162443_1e097c79_8958a65f
0e_7a6d9b0b__00000000_95aefe44_693868f3_ae445cca_b093df3b_e4c5244e_9f459a20_8d8d5c0b_b7fc7fc0_0683ab57_33a4289e_ee7ca9a7_fbd237fa_2a7b62da_7a6d9b0b_05fb991e_76f15d5d_974251c3_a22c7cf8_6282990b_50f6b395_4d24c9a9_378472ee_e66ba7c1_46e91766_0d056ce8_c72cb5ab_00000000_00000000_4b162443_1e097c79_8958a65f
1d_63d2a87f__00000000_95aefe44_693868f3_ae445cca_b093df3b_e4c5244e_9f459a20_8d8d5c0b_b7fc7fc0_0683ab57_33a4289e_ee7ca9a7_fbd237fa_2a7b62da_7a6d9b0b_05fb991e_76f15d5d_974251c3_a22c7cf8_6282990b_50f6b395_4d24c9a9_378472ee_e66ba7c1_46e91766_0d056ce8_c72cb5ab_00000000_00000000_63d2a87f_1e097c79_8958a65f
1f_6c4ecfd6__00000000_95aefe44_693868f3_ae445cca_b093df3b_e4c5244e_9f459a20_8d8d5c0b_b7fc7fc0_0683ab57_33a4289e_ee7ca9a7_fbd237fa_2a7b62da_7a6d9b0b_05fb991e_76f15d5d_974251c3_a22c7cf8_6282990b_50f6b395_4d24c9a9_378472ee_e66ba7c1_46e91766_0d056ce8_c72cb5ab_00000000_00000000_63d2a87f_1e097c79_6c4ecfd6
0d_82028106__00000000_95aefe44_693868f3_ae445cca_b093df3b_e4c5244e_9f459a20_8d8d5c0b_b7fc7fc0_0683ab57_33a4289e_ee7ca9a7_fbd237fa_82028106_7a6d9b0b_05fb991e_76f15d5d_974251c3_a22c7cf8_6282990b_50f6b395_4d24c9a9_378472ee_e66ba7c1_46e91766_0d056ce8_c72cb5ab_00000000_00000000_63d2a87f_1e097c79_6c4ecfd6
11_29e08cf4__00000000_95aefe44_693868f3_ae445cca_b093df3b_e4c5244e_9f459a20_8d8d5c0b_b7fc7fc0_0683ab57_33a4289e_ee7ca9a7_fbd237fa_82028106_7a6d9b0b_05fb991e_76f15d5d_29e08cf4_a22c7cf8_6282990b_50f6b395_4d24c9a9_378472ee_e66ba7c1_46e91766_0d056ce8_c72cb5ab_00000000_00000000_63d2a87f_1e097c79_6c4ecfd6
01_93b508e7__00000000_93b508e7_693868f3_ae445cca_b093df3b_e4c5244e_9f459a20_8d8d5c0b_b7fc7fc0_0683ab57_33a4289e_ee7ca9a7_fbd237fa_82028106_7a6d9b0b_05fb991e_76f15d5d_29e08cf4_a22c7cf8_6282990b_50f6b395_4d24c9a9_378472ee_e66ba7c1_46e91766_0d056ce8_c72cb5ab_00000000_00000000_63d2a87f_1e097c79_6c4ecfd6
14_082d866c__00000000_93b508e7_693868f3_ae445cca_b093df3b_e4c5244e_9f459a20_8d8d5c0b_b7fc7fc0_0683ab57_33a4289e_ee7ca9a7_fbd237fa_82028106_7a6d9b0b_05fb991e_76f15d5d_29e08cf4_a22c7cf8_6282990b_082d866c_4d24c9a9_378472ee_e66ba7c1_46e91766_0d056ce8_c72cb5ab_00000000_00000000_63d2a87f_1e097c79_6c4ecfd6
12_b98cc6c0__00000000_93b508e7_693868f3_ae445cca_b093df3b_e4c5244e_9f459a20_8d8d5c0b_b7fc7fc0_0683ab57_33a4289e_ee7ca9a7_fbd237fa_82028106_7a6d9b0b_05fb991e_76f15d5d_29e08cf4_b98cc6c0_6282990b_082d866c_4d24c9a9_378472ee_e66ba7c1_46e91766_0d056ce8_c72cb5ab_00000000_00000000_63d2a87f_1e097c79_6c4ecfd6
08_b112b2eb__00000000_93b508e7_693868f3_ae445cca_b093df3b_e4c5244e_9f459a20_8d8d5c0b_b112b2eb_0683ab57_33a4289e_ee7ca9a7_fbd237fa_82028106_7a6d9b0b_05fb991e_76f15d5d_29e08cf4_b98cc6c0_6282990b_082d866c_4d24c9a9_378472ee_e66ba7c1_46e91766_0d056ce8_c72cb5ab_00000000_00000000_63d2a87f_1e097c79_6c4ecfd6
1a_beda90bd__00000000_93b508e7_693868f3_ae445cca_b093df3b_e4c5244e_9f459a20_8d8d5c0b_b112b2eb_0683ab57_33a4289e_ee7ca9a7_fbd237fa_82028106_7a6d9b0b_05fb991e_76f15d5d_29e08cf4_b98cc6c0_6282990b_082d866c_4d24c9a9_378472ee_e66ba7c1_46e91766_0d056ce8_beda90bd_00000000_00000000_63d2a87f_1e097c79_6c4ecfd6
0b_34c2bf43__00000000_93b508e7_693868f3_ae445cca_b093df3b_e4c5244e_9f459a20_8d8d5c0b_b112b2eb_0683ab57_33a4289e_34c2bf43_fbd237fa_82028106_7a6d9b0b_05fb991e_76f15d5d_29e08cf4_b98cc6c0_6282990b_082d866c_4d24c9a9_378472ee_e66ba7c1_46e91766_0d056ce8_beda90bd_00000000_00000000_63d2a87f_1e097c79_6c4ecfd6
05_d09de25a__00000000_93b508e7_693868f3_ae445cca_b093df3b_d09de25a_9f459a20_8d8d5c0b_b112b2eb_0683ab57_33a4289e_34c2bf43_fbd237fa_82028106_7a6d9b0b_05fb991e_76f15d5d_29e08cf4_b98cc6c0_6282990b_082d866c_4d24c9a9_378472ee_e66ba7c1_46e91766_0d056ce8_beda90bd_00000000_00000000_63d2a87f_1e097c79_6c4ecfd6
0b_410ded3b__00000000_93b508e7_693868f3_ae445cca_b093df3b_d09de25a_9f459a20_8d8d5c0b_b112b2eb_0683ab57_33a4289e_410ded3b_fbd237fa_82028106_7a6d9b0b_05fb991e_76f15d5d_29e08cf4_b98cc6c0_6282990b_082d866c_4d24c9a9_378472ee_e66ba7c1_46e91766_0d056ce8_beda90bd_00000000_00000000_63d2a87f_1e097c79_6c4ecfd6
0a_6d0360e0__00000000_93b508e7_693868f3_ae445cca_b093df3b_d09de25a_9f459a20_8d8d5c0b_b112b2eb_0683ab57_6d0360e0_410ded3b_fbd237fa_82028106_7a6d9b0b_05fb991e_76f15d5d_29e08cf4_b98cc6c0_6282990b_082d866c_4d24c9a9_378472ee_e66ba7c1_46e91766_0d056ce8_beda90bd_00000000_00000000_63d2a87f_1e097c79_6c4ecfd6
0f_380440a4__00000000_93b508e7_693868f3_ae445cca_b093df3b_d09de25a_9f459a20_8d8d5c0b_b112b2eb_0683ab57_6d0360e0_410ded3b_fbd237fa_82028106_7a6d9b0b_380440a4_76f15d5d_29e08cf4_b98cc6c0_6282990b_082d866c_4d24c9a9_378472ee_e66ba7c1_46e91766_0d056ce8_beda90bd_00000000_00000000_63d2a87f_1e097c79_6c4ecfd6
1f_6e31fef2__00000000_93b508e7_693868f3_ae445cca_b093df3b_d09de25a_9f459a20_8d8d5c0b_b112b2eb_0683ab57_6d0360e0_410ded3b_fbd237fa_82028106_7a6d9b0b_380440a4_76f15d5d_29e08cf4_b98cc6c0_6282990b_082d866c_4d24c9a9_378472ee_e66ba7c1_46e91766_0d056ce8_beda90bd_00000000_00000000_63d2a87f_1e097c79_6e31fef2
04_fd0ca385__00000000_93b508e7_693868f3_ae445cca_fd0ca385_d09de25a_9f459a20_8d8d5c0b_b112b2eb_0683ab57_6d0360e0_410ded3b_fbd237fa_82028106_7a6d9b0b_380440a4_76f15d5d_29e08cf4_b98cc6c0_6282990b_082d866c_4d24c9a9_378472ee_e66ba7c1_46e91766_0d056ce8_beda90bd_00000000_00000000_63d2a87f_1e097c79_6e31fef2
1b_10b39ac1__00000000_93b508e7_693868f3_ae445cca_fd0ca385_d09de25a_9f459a20_8d8d5c0b_b112b2eb_0683ab57_6d0360e0_410ded3b_fbd237fa_82028106_7a6d9b0b_380440a4_76f15d5d_29e08cf4_b98cc6c0_6282990b_082d866c_4d24c9a9_378472ee_e66ba7c1_46e91766_0d056ce8_beda90bd_10b39ac1_00000000_63d2a87f_1e097c79_6e31fef2
0a_58befbc4__00000000_93b508e7_693868f3_ae445cca_fd0ca385_d09de25a_9f459a20_8d8d5c0b_b112b2eb_0683ab57_58befbc4_410ded3b_fbd237fa_82028106_7a6d9b0b_380440a4_76f15d5d_29e08cf4_b98cc6c0_6282990b_082d866c_4d24c9a9_378472ee_e66ba7c1_46e91766_0d056ce8_beda90bd_10b39ac1_00000000_63d2a87f_1e097c79_6e31fef2
0a_298e7114__00000000_93b508e7_693868f3_ae445cca_fd0ca385_d09de25a_9f459a20_8d8d5c0b_b112b2eb_0683ab57_298e7114_410ded3b_fbd237fa_82028106_7a6d9b0b_380440a4_76f15d5d_29e08cf4_b98cc6c0_6282990b_082d866c_4d24c9a9_378472ee_e66ba7c1_46e91766_0d056ce8_beda90bd_10b39ac1_00000000_63d2a87f_1e097c79_6e31fef2
18_df55c596__00000000_93b508e7_693868f3_ae445cca_fd0ca385_d09de25a_9f459a20_8d8d5c0b_b112b2eb_0683ab57_298e7114_410ded3b_fbd237fa_82028106_7a6d9b0b_380440a4_76f15d5d_29e08cf4_b98cc6c0_6282990b_082d866c_4d24c9a9_378472ee_e66ba7c1_df55c596_0d056ce8_beda90bd_10b39ac1_00000000_63d2a87f_1e097c79_6e31fef2
10_bf618501__00000000_93b508e7_693868f3_ae445cca_fd0ca385_d09de25a_9f459a20_8d8d5c0b_b112b2eb_0683ab57_298e7114_410ded3b_fbd237fa_82028106_7a6d9b0b_380440a4_bf618501_29e08cf4_b98cc6c0_6282990b_082d866c_4d24c9a9_378472ee_e66ba7c1_df55c596_0d056ce8_beda90bd_10b39ac1_00000000_63d2a87f_1e097c79_6e31fef2
0d_4d848450__00000000_93b508e7_693868f3_ae445cca_fd0ca385_d09de25a_9f459a20_8d8d5c0b_b112b2eb_0683ab57_298e7114_410ded3b_fbd237fa_4d848450_7a6d9b0b_380440a4_bf618501_29e08cf4_b98cc6c0_6282990b_082d866c_4d24c9a9_378472ee_e66ba7c1_df55c596_0d056ce8_beda90bd_10b39ac1_00000000_63d2a87f_1e097c79_6e31fef2
01_f15c8f6f__00000000_f15c8f6f_693868f3_ae445cca_fd0ca385_d09de25a_9f459a20_8d8d5c0b_b112b2eb_0683ab57_298e7114_410ded3b_fbd237fa_4d848450_7a6d9b0b_380440a4_bf618501_29e08cf4_b98cc6c0_6282990b_082d866c_4d24c9a9_378472ee_e66ba7c1_df55c596_0d056ce8_beda90bd_10b39ac1_00000000_63d2a87f_1e097c79_6e31fef2
00_c9d61f75__00000000_f15c8f6f_693868f3_ae445cca_fd0ca385_d09de25a_9f459a20_8d8d5c0b_b112b2eb_0683ab57_298e7114_410ded3b_fbd237fa_4d848450_7a6d9b0b_380440a4_bf618501_29e08cf4_b98cc6c0_6282990b_082d866c_4d24c9a9_378472ee_e66ba7c1_df55c596_0d056ce8_beda90bd_10b39ac1_00000000_63d2a87f_1e097c79_6e31fef2
12_d095c032__00000000_f15c8f6f_693868f3_ae445cca_fd0ca385_d09de25a_9f459a20_8d8d5c0b_b112b2eb_0683ab57_298e7114_410ded3b_fbd237fa_4d848450_7a6d9b0b_380440a4_bf618501_29e08cf4_d095c032_6282990b_082d866c_4d24c9a9_378472ee_e66ba7c1_df55c596_0d056ce8_beda90bd_10b39ac1_00000000_63d2a87f_1e097c79_6e31fef2
